------------------------------------- 

--KTU 2015

--Informatikos fakultetas
--Kompiuteriu katedra
--Kompiuteriu Architektura [P175B125] 
--Kazimieras Bagdonas 

--v1.0

------------------------------------- 
--KTU 2016 

--ditto

--v1.01
--panaikinta "save" mikrokomanda registrams, sutrumpinta ROM eilute nuo 75 iki 69 bitu, nesuderinama su V1.0   

------------------------------------- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
	port (
		RST_ROM : in std_logic;
		ROM_CMD : in std_logic_vector(7 downto 0);  
		ROM_Dout : out std_logic_vector(1 to 69)
		);
end ROM ;

architecture rtl of ROM is
	
	type memory is array (0 to 255) of std_logic_vector(1 to 69) ; 
	
	constant ROM_CMDln : memory := (  
--                    1         2         3         4         5         6            Dvi komentaro eilutes duoda bitu numerius   
--           123456789012345678901234567890123456789012345678901234567890123456789    (nuo 1 iki 69)
0=> "010000000000000100000000000000000000000000000000000000000000000000000",  --B = N1
1=> "010000000000000000000010000000000000000000000000000000000000000000000",  --C = N2
2=> "000010000000000000000000000000000000000000000000000000000000000000000",  --MUX = C
3=> "000000001000000000000000000000000000000000000000000100000000000000000",  --M = not L, A = M
4=> "001000000000000000000010000001000000000000000000000000000000000000000",  --MUX = A, C = A, D = A
5=> "000000000000000000000000000000000000000000000000000000000010000000000",  --RESET(A)
6=> "000010000000000000000000000000000000000000000000000000000000000000000",  --MUX = C
7=> "110000000100100000000000000000000000000000000000000000000000000000000",  --LS = 8
8=> "000000001000000000000000000000000000000000000000001000000000000000000",  --M = L + R, A = M
9=> "000000000000000000000000000000000000000000000000000000000000000000001",  --CNT--
10=> "000000000000000000000001000000010000000000000000000000000000000000000",  --LL1(C), LR1(D)
11=> "111010000011100000000000000000000000000000000000000000000000000000000",  --LS = 13
12=> "001000000000000000000000000000000000000000000000000000000000000000000",  --MUX = A
13=> "000000001000000000000000000000000000000000000000000100000000000000000",  --M = not L, A = M
14=> "000100000000000000000000000000000000000000000000000000000000000000000",  --MUX = B
15=> "000000001000000000000000000000000000000000000000001000000000000000000",  --M = L + R, A = M
16=> "001000000000000000000000000000000000000000000000000000000000000000000",  --MUX = A
17=> "000000000000000000000000000000000000000000000000000000000000000000010",  --DOUT









	
	others => (others => '0') );   
	
	
	
begin
	process (RST_ROM, ROM_CMD) 
		
	begin
		if RST_ROM'event and RST_ROM = '1' then 
			ROM_Dout <= ROM_CMDln(0);
		elsif ROM_CMD'event then
			ROM_Dout <= ROM_CMDln(to_integer(unsigned(ROM_CMD))); 
		end if;
		
	end process;
	
end rtl;